package rf_agent_pkg;

  //uvm pakage and macros
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  


`include "rf_item.sv"
`include "rf_agent_cfg.sv"
`include "rf_monitor.sv"
`include "rf_driver.sv"
`include "rf_reg2hmc_adapter.sv"
`include "rf_sequencer.sv"
`include "rf_agent.sv"


endpackage : rf_agent_pkg