//`include "axi_interface.sv"

package axi_pkg;
`include "uvm_macros.svh"
import uvm_pkg::*;
import cmd_pkg::*;

`include "axi_config.svh"
`include "valid_data.svh"
`include "hmc_pkt_item_request.svh"
`include "axi_sequencer.svh"
`include "axi_driver.svh"
`include "axi_monitor.svh"
`include "axi_agent.svh" 


endpackage : axi_pkg
