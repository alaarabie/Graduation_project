package rf_reg_block_pkg;
  
  //uvm pakage and macros
  import uvm_pkg::*;
  `include "uvm_macros.svh"


`include "reg_error_abort_not_cleared.svh"
`include "reg_counter_reset.svh"
`include "reg_errors_on_rx.svh"
`include "reg_poisoned_packets.svh"
`include "reg_rcvd_rsp.svh"
`include "reg_run_length_bit_flip.svh"
`include "reg_sent_np.svh"
`include "reg_sent_p.svh"
`include "reg_sent_r.svh"
`include "reg_status_general.svh"
`include "reg_status_init.svh"
`include "reg_tx_link_retries.svh"
`include "reg_control.svh"

`include "rf_reg_block.svh"
  
endpackage : rf_reg_block_pkg