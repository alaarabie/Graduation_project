package test_pkg ;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
    import cmd_pkg::*;
    import tb_pkg::* ;

	`include "vseq_base.sv"
	`include "hmc_vseq.sv"
	`include "base_test.sv"
	`include "random_test.sv"	


endpackage : test_pkg