package seq_pkg ;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
    import cmd_pkg::*;
    import axi_pkg::* ;    
    import hmc_agent_pkg::* ;
    import rf_reg_block_pkg::* ;    
    import rf_agent_pkg::* ;
    // import test_pkg::* ;
    import tb_pkg::* ;


    `include "base_seq.sv"
    `include "hmc_initialization_seq.sv"    
    `include "hmc_response_seq.sv"            
    `include "hmc_state_seq.sv" 
    `include "rf_control_configuration_seq.sv"
    `include "rf_control_read_seq.sv"
    `include "rf_counters_seq.sv"
    `include "rf_status_general_seq.sv"
    `include "rf_control_sleep_seq.sv" 
    `include "rf_reset_seq.sv" 
    `include "rf_status_init_mirror_seq.sv"            
    `include "axi_seq.sv"   
   

endpackage : seq_pkg