package tb_pkg ;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
    import cmd_pkg::*;
    import axi_pkg::* ;
    import hmc_agent_pkg::* ;
    import rf_reg_block_pkg::* ;    
    import rf_agent_pkg::* ;
    import tb_params_pkg::* ;

  `include "coverage.svh"
  `include "scoreboard.svh"
	`include "env_cfg.svh"
	`include "vsequencer.svh"	
	`include "env.svh"    

endpackage : tb_pkg