interface hmc_agent_if



endinterface : hmc_agent_if