interface system_if (input clk);

logic           res_n;    //output

endinterface : system_if