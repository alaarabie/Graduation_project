package seq_pkg ;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
    import cmd_pkg::*;
    import axi_pkg::* ;    
    import hmc_agent_pkg::* ;
    import rf_reg_block_pkg::* ;    
    import rf_agent_pkg::* ;
    import tb_pkg::* ;


    `include "base_seq.svh"  
           
    `include "rf_control_read_seq.svh"
    `include "rf_counters_seq.svh"
    `include "rf_status_general_seq.svh"
    `include "rf_control_sleep_seq.svh" 
    `include "rf_status_init_seq.svh"
    `include "initialization_seq.svh"
    `include "rf_wrong_op_seq.svh"
                 
    `include "axi_base_seq.svh" 
    `include "axi_read_seq.svh"  
    `include "axi_posted_seq.svh" 
    `include "axi_write_seq.svh" 

    `include "reset-sequences/reset1_seq.svh" 
    `include "reset-sequences/reset2_seq.svh" 
    `include "reset-sequences/reset3_seq.svh" 
    `include "reset-sequences/reset4_seq.svh" 
    `include "reset-sequences/reset5_seq.svh" 
   

endpackage : seq_pkg