package rf_agent_pkg;

  //uvm pakage and macros
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  


`include "rf_item.svh"
`include "rf_agent_cfg.svh"
`include "rf_monitor.svh"
`include "rf_driver.svh"
`include "rf_reg2openhmc_adapter.svh"
`include "rf_sequencer.svh"
`include "rf_agent.svh"


endpackage : rf_agent_pkg