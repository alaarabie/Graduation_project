package tb_pkg ;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
    import cmd_pkg::*;
    import axi_pkg::* ;
    import hmc_agent_pkg::* ;
    import rf_reg_block_pkg::* ;    
    import rf_agent_pkg::* ;
    import tb_params_pkg::* ;

    
	`include "env_cfg.sv"
	`include "vsequencer.sv"	
	`include "env.sv"    

    // import seq_pkg::* ;
    // import test_pkg::* ;

endpackage : tb_pkg